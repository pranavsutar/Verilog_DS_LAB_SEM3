//written by Mathew K J CS20B021

module ANDgate_2in(A,B,C);

input A;
input B;

output C;

assign C = A&B;

endmodule //ANDgate_2in