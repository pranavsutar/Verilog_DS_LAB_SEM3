// Written BY CS20BO29

module ANDgate_2_inputs (a,b,y);

input a;
imput b;

output y;

assign y = a & b;

endmodule